// module arbiter(
//     input wire clock,
//     input wire reset,

//     input
// );

// endmodule